package comp_cic_tsb_pkg; 
 
integer test_case = 2; // #case for test 
 
parameter Win = 16; 
parameter Wcoef = 18; 
parameter Wout = 34; 
parameter Ng = 18; 
parameter Num_coef = 17; 
 
endpackage