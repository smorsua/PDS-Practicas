package cic_tsb_pkg; 
 
integer test_case = 3; // #case for test 
 
parameter Win = 18; 
parameter Ncomb = 1; 
parameter Ng = 27; 
parameter Wout = 48; 
parameter R = 2000; 
 
endpackage