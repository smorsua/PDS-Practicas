package cic_tsb_pkg; 
 
integer test_case = 1; // #case for test 
 
parameter Win = 18; 
parameter Ncomb = 1; 
parameter Ng = 27; 
parameter Wout = 16; 
parameter R = 2000; 
 
endpackage