package dp_mod_tsb_pkg; 
 
integer test_case = 1; // #case for test 
integer in_sample_num = 38401; // #processed input samples 
 
integer fsc = 96; // Clock frequency (MHz) 
integer fmod = 5; // Modulation frequency (kHz) 
integer fc = 1.070000e+01; // Carrier frequency (MHz) 
integer im_am = 32767; // AM modulation index 
integer im_fm = 0; // FM modulation index (not used in AM) 
 
endpackage