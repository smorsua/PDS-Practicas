package dp_mod_tsb_pkg; 
 
integer test_case = 2; // #case for test 
integer in_sample_num = 19201; // #processed input samples 
 
integer fsc = 96; // Clock frequency (MHz) 
integer fmod = 5; // Modulation frequency (kHz) 
integer fc = 1; // Carrier frequency (MHz) 
integer im_am = 0; // AM modulation index (not used in FM) 
integer im_fm = 478; // FM modulation index (kHz) 
 
endpackage